// --------------------------------------------------------------------
//
// --------------------------------------------------------------------

module bit_serial_adder
( input  clk
, input  reset
, input  a
, input  b
, output x
);
  // --------------------------------------------------------------------
  wire c_in;
  wire sum;
  wire c_out;

  full_adder fa_i(.*);

  // --------------------------------------------------------------------
  d_flip_flop ff_c_in_i(.d(c_out), .q(c_in), .q_n(), .*);
  d_flip_flop ff_sum_i (.d(sum)  , .q(x)   , .q_n(), .*);

// --------------------------------------------------------------------
endmodule
