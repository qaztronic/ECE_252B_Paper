// --------------------------------------------------------------------
//
// --------------------------------------------------------------------

package tb_top_pkg;

  // --------------------------------------------------------------------
  function void test_done(string test_pass);
    $display("--------------------------------------------------------------------");
    $display("Test %s!!!", test_pass);
    $stop;
  endfunction

// --------------------------------------------------------------------
endpackage

