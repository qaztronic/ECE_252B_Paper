// --------------------------------------------------------------------
//
// --------------------------------------------------------------------

module d_flip_flop
( input  clk
, input  d
, input  reset
, output reg q
, output q_n
);
  // --------------------------------------------------------------------
  assign q_n = ~q;

  always_ff @(posedge clk)
    if(reset)
      q <= 0;
    else
      q <= d;

// --------------------------------------------------------------------
endmodule
