// --------------------------------------------------------------------
//
// --------------------------------------------------------------------

module counter_5_to_3
( input [4:1] x
, input c_in
, output s
, output c
, output c_out
);
  // --------------------------------------------------------------------
  wire x_lo = x[1] ^ x[2];
  wire x_hi = x[3] ^ x[4];
  wire x_all = x_lo ^ x_hi;
  
  // --------------------------------------------------------------------
  // m0(in0, in1, sel, out);
  
  // --------------------------------------------------------------------
  wire m0_out;
  mux m0(x[1], x[3], x_lo, m0_out);

  // --------------------------------------------------------------------
  wire m1_out;
  mux m1(x[4], c_in, x_all, m1_out);

  
  // --------------------------------------------------------------------
  assign c_out = m0_out;
  assign s = x_all ^ c_in;
  assign c = m1_out;
  
  
  // // --------------------------------------------------------------------
  // wire 
  
  // full_adder fa0
  // ( .a    (x[0])
  // , .b    (x[1])
  // , .c_in (x[2])
  // , .sum  ()
  // , .c_out()
  // );
  
  // // --------------------------------------------------------------------
  // full_adder fa1
  // ( input  a
  // , input  b
  // , input  c_in
  // , output sum
  // , output c_out
  // );
  
  // // --------------------------------------------------------------------
  // full_adder fa1
  // ( input  a
  // , input  b
  // , input  c_in
  // , output sum
  // , output c_out
  // );
  
  
  // // --------------------------------------------------------------------
  // // m0(in0, in1, sel, out);
  // wire m0_out;
  // mux m0(x[4], ~x[4], x[3], m0_out);

  // // --------------------------------------------------------------------
  // wire m1_out;
  // mux m1(x[2], ~x[2], x[1], m1_out);

  // // --------------------------------------------------------------------
  // wire m2_out = m0_out;
  // // mux m2(in0, in1, sel, m2_out);

  // // --------------------------------------------------------------------
  // wire m3_out;
  // mux m3(x[1], x[3], m1_out, m3_out);

  // // --------------------------------------------------------------------
  // wire m4_out;
  // mux m4(x[4], c_in, m2_out, m4_out);

  // // --------------------------------------------------------------------
  // wire m5_out;
  // mux m5(c_in, ~c_in, m2_out, m5_out);

  // // --------------------------------------------------------------------
  // // assign sum   = {m4_out, m5_out};
  // assign c_out = m3_out;
  // assign s = m5_out;
  // assign c = m4_out;

// --------------------------------------------------------------------
endmodule
