// --------------------------------------------------------------------
//
// --------------------------------------------------------------------

module cell #(N, W)
( input  clk
, input  reset
, input  left_in
, input  right_in
, input  top_in
, input  bottom_in
, output left_out
, output right_out
, output top_out
, output bottom_out
);
  // --------------------------------------------------------------------
  import alu_pkg::*;
  
  // --------------------------------------------------------------------

// --------------------------------------------------------------------
endmodule

