// --------------------------------------------------------------------
//
// --------------------------------------------------------------------

module counter_5_to_3
( input [4:1] x
, input c_in
, output s
, output c
, output c_out
);
  // --------------------------------------------------------------------
  wire hi_sum;
  wire hi_c_out;

  full_adder fa_hi
  ( .a    (x[3])
  , .b    (x[4])
  , .c_in (c_in)
  , .sum  (hi_sum)
  , .c_out(hi_c_out)
  );

  // --------------------------------------------------------------------
  wire lo_c_out;

  full_adder fa_lo
  ( .a    (x[1])
  , .b    (x[2])
  , .c_in (hi_sum)
  , .sum  (s)
  , .c_out(lo_c_out)
  );

  // --------------------------------------------------------------------
  assign c_out = hi_c_out & lo_c_out; // half adder
  assign c = hi_c_out ^ lo_c_out;

// --------------------------------------------------------------------
endmodule
