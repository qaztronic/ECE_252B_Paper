// --------------------------------------------------------------------
//
// --------------------------------------------------------------------

package alu_pkg;

  // --------------------------------------------------------------------

  enum logic [3:0]
    {
      GET_WORD_IN   = 3'b001,
      MUX_WORD_OUT  = 3'b010,
      LAST_WORD_OUT = 3'b100
    } alu_op;

// --------------------------------------------------------------------
endpackage

